package eportrxdrv_pkg;

    `include "classes.sv"

endpackage
